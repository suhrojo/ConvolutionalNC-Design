`default_nettype none

module FCL ( // Full Connected Layer
    input wire [7:0] data_in,
    input wire clk,
    input wire rst_n, 

    output reg [7:0] data_out
);

endmodule