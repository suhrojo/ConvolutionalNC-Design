`default_nettype none

module PoolingLayer(
input wire clk,
input wire rst_n,
input wire [7:0] data_in

output wire [7:0] data_out
);

endmodule;