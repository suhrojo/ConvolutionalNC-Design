`default_nettype 

module HiddenLayer(

);

endmodule